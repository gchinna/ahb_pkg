`ifndef _AHP_MACROS_SVH 
`define _AHP_MACROS_SVH 

  `ifndef AHB_AWIDTH
    `define AHB_AWIDTH 32  // default addr width
  `endif

  `ifndef AHB_DWIDTH
    `define AHB_DWIDTH 32  // default data width
  `endif

 
`endif // _AHP_MACROS_SVH
